-- very simple tb to create an input packets to the slave port

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
USE ieee.numeric_std.ALL; 

entity tb is
end tb;

architecture tb of tb is
    -- change here if you want to send longer packets
    constant MAX_FLITS : integer := 4;

	signal clock:    std_logic := '0';
	signal reset:    std_logic;  

	-- axi slave streaming interface
	signal s_valid_i :  std_logic;
	signal s_ready_o :  std_logic;
	signal s_last_i  :  std_logic;
	signal s_data_i  :  std_logic_vector(31 downto 0);

	-- axi master streaming interface
	signal m_valid_o :  std_logic;
	signal m_ready_i :  std_logic;
	signal m_last_o  :  std_logic;
	signal m_data_o  :  std_logic_vector(31 downto 0);
           

    type packet_t is array (0 to MAX_FLITS+1) of std_logic_vector(31 downto 0);	
	
	-- send one work according to the AXI Streaming master protocol
	procedure SendFlit(signal clock  : in  std_logic;
	                   constant flit : in  std_logic_vector(31 downto 0);
	                   --- AXI master streaming 
	                   signal data   : out std_logic_vector(31 downto 0);
	                   signal valid  : out std_logic;
	                   signal last   : out std_logic;
	                   constant end_of_packet   : in std_logic;
	                   signal ready  : in  std_logic
	                   ) is
	begin
		wait until rising_edge(clock);
		-- If both the AXI interface and the router runs at the rising edge, then it is necessary to add 
		--   a delay at the inputs. The solution was to put an inverted in the clock in the Router_Board entity. 
		-- This way the delay is not necessary and it is also not necessary to change the router's vhdl   
        data <= flit;
        valid <= '1';
        last <= end_of_packet;
        wait for 8ns; -- simulate delay at the primary inputs
        while ready /= '1' loop
             wait until falling_edge(clock); -- data is buffered at the falling edge
        end loop;	
	end procedure;
	
	procedure SendPacket(signal clock  : in  std_logic;
                       constant packet : in  packet_t;
                       --- AXI master streaming 
                       signal data   : out std_logic_vector(31 downto 0);
                       signal valid  : out std_logic;
                       signal last   : out std_logic;
                       signal ready  : in  std_logic
                       ) is
        variable num_flits : integer;
    begin
         -- send header
        SendFlit(clock,packet(0),data,valid,last,'0',ready);
        -- send size
        SendFlit(clock,packet(1),data,valid,last,'0',ready);
        num_flits := to_integer(signed(packet(1)));
        -- send payload
        for f in 2 to num_flits loop
            SendFlit(clock,packet(f),data,valid,last,'0',ready);
        end loop;
        SendFlit(clock,packet(num_flits+1),data,valid,last,'1',ready);
        
      -- end of the packet transfer
        wait until rising_edge(clock);
        wait for 4 ns;
        last <= '0';
        valid <= '0';
        data <= (others => '0');
        -- wait a while to start the next packet transfer 
        wait for 100 ns;    
    end procedure;

	
begin

	reset <= '0', '1' after 100 ns; -- active low

    -- 50 MHz, as the default freq generated by the PS
	process
	begin
		clock <= not clock;
		wait for 10 ns;
		clock <= not clock;
		wait for 10 ns;
	end process;
	
	-- the master ports is always ready to receive
	m_ready_i <= '1';

    ----------------------------------------------------
    -- send packets to the slave port
    ----------------------------------------------------
    process
         variable  packet : packet_t;
	begin
	    s_valid_i <= '0';
		s_data_i <= (others => '0');
		s_last_i <= '0';
		wait for 200 ns;
		wait until rising_edge(clock);
		
		-- from the east to local
		packet := (x"00000101", x"00000002", x"00000000", x"00000001", x"00000000", x"00000000");
		SendPacket(clock, packet, s_data_i, s_valid_i, s_last_i, s_ready_o);
		-- from the north to local
        packet := (x"00000101", x"00000002", x"00000001", x"00000002", x"00000000", x"00000000");
        SendPacket(clock, packet, s_data_i, s_valid_i, s_last_i, s_ready_o);
		-- from the west to local
        packet := (x"00000101", x"00000004", x"00000000", x"11111111", x"22222222", x"33333333");
        SendPacket(clock, packet, s_data_i, s_valid_i, s_last_i, s_ready_o);
		-- from the south to local
        packet := (x"00000101", x"00000004", x"00000001", x"44444444", x"55555555", x"66666666");
        SendPacket(clock, packet, s_data_i, s_valid_i, s_last_i, s_ready_o);
		
		-- block here. do not send it again
		wait;
	end process;


 router: entity work.noc_counter
  port map ( 
        clock     => clock,
        reset_n   => reset,
	-- axi slave streaming interface
        s_valid_i => s_valid_i,
        s_ready_o => s_ready_o,
        s_last_i  => s_last_i,
        s_data_i  => s_data_i,
        -- axi master streaming interface
        m_valid_o => m_valid_o,
        m_ready_i => m_ready_i,
        m_last_o  => m_last_o,
        m_data_o  => m_data_o
	);
	
end tb;

